library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity lab3 is
  port(CLOCK_50            : in  std_logic;
       KEY                 : in  std_logic_vector(3 downto 0);
       SW                  : in  std_logic_vector(17 downto 0);
       VGA_R, VGA_G, VGA_B : out std_logic_vector(9 downto 0);  -- The outs go to VGA controller
       VGA_HS              : out std_logic;
       VGA_VS              : out std_logic;
       VGA_BLANK           : out std_logic;
       VGA_SYNC            : out std_logic;
       VGA_CLK             : out std_logic);
end lab3;

architecture rtl of lab3 is

 --Component from the Verilog file: vga_adapter.v

  component vga_adapter
    generic(RESOLUTION : string);
    port (resetn                                       : in  std_logic;
          clock                                        : in  std_logic;
          colour                                       : in  std_logic_vector(2 downto 0);
          x                                            : in  std_logic_vector(7 downto 0);
          y                                            : in  std_logic_vector(6 downto 0);
          plot                                         : in  std_logic;
          VGA_R, VGA_G, VGA_B                          : out std_logic_vector(9 downto 0);
          VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_CLK : out std_logic);
  end component;

  signal x      : std_logic_vector(7 downto 0);
  signal y      : std_logic_vector(6 downto 0);
  signal colour : std_logic_vector(2 downto 0);
  signal plot   : std_logic;

  signal clock, reset_async : std_logic;

begin
  
  clock       <= clock_50;
  reset_async <= not key(3);
  plot   <= not KEY(0);

  -- includes the vga adapter, which should be in your project 

  vga_u0 : vga_adapter
    generic map(RESOLUTION => "160x120") 
    port map(resetn    => KEY(3),
             clock     => CLOCK_50,
             colour    => colour,
             x         => x,
             y         => y,
             plot      => plot,
             VGA_R     => VGA_R,
             VGA_G     => VGA_G,
             VGA_B     => VGA_B,
             VGA_HS    => VGA_HS,
             VGA_VS    => VGA_VS,
             VGA_BLANK => VGA_BLANK,
             VGA_SYNC  => VGA_SYNC,
             VGA_CLK   => VGA_CLK);

    process(clock, reset_async)
    variable x_count : unsigned(7 downto 0) := "00000000";
    variable y_count : unsigned(6 downto 0) := "0000000";
    begin
      x <= std_logic_vector(x_count);
      y <= std_logic_vector(y_count);
      if (rising_edge(clock)) then
        y_count := y_count + 1;
        if (y_count mod 120 = 0) then
          y_count := "0000000";
          x_count := x_count + 1;
        end if;
        if (x_count mod 160 = 0) then
          x_count := "00000000";
        end if;
        if (reset_async = '1') then
          x_count := "00000000";
          y_count := "0000000";
        end if;
        case (y_count mod 8) is
          when "0000000" => colour <= "001";
          when "0000001" => colour <= "010";
          when "0000010" => colour <= "011";
          when "0000011" => colour <= "100";
          when "0000100" => colour <= "101";
          when "0000101" => colour <= "110";
          when "0000110" => colour <= "111";
          when "0000111" => colour <= "000";
          when others => colour <= "000";
        end case;
      end if;
    end process;
end rtl;


